-- State Machine

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY StateMachine IS
	PORT( CLK, BUTTON, REG_9, REG_0, COUNT: IN STD_LOGIC;
			SL, SR: OUT STD_LOGIC);
END StateMachine;

ARCHITECTURE rtl OF StateMachine IS

	TYPE state IS (INIT, ShiftLeft, ShiftRight);
	SIGNAL current_state: state := INIT;
	SIGNAL next_state: state;
	
	
BEGIN

	PROCESS(CLK)
	BEGIN
		IF (CLK' EVENT) AND (CLK = '1') THEN
			CASE current_state IS
				WHEN INIT =>
					SL <= '0';
					SR <= '0';
					IF BUTTON = '0' THEN
						next_state <= INIT;
					ELSE 
						next_state <= ShiftLeft;
					END IF;
					
				WHEN ShiftLeft =>
					SL <= '1';
					SR <= '0';
					IF REG_9 = '1' THEN
						next_state <= ShiftRight;
					ELSE 
						next_state <= ShiftLeft;
					END IF;
					
				WHEN ShiftRight =>
					SL <= '0';
					SR <= '1';
					IF REG_0 = '1' THEN
						next_state <= ShiftLeft;
					ELSE 
						next_state <= ShiftRight;
					END IF;
			END CASE;
		END IF;
	END PROCESS;
END rtl;
		