-- Counter

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Counter IS
	PORT( CLK, ASYNCCLRN, SYNCCLRN : IN STD_LOGIC;
			Q : OUT STD_LOGIC_VECTOR(19 DOWNTO 0));
END Counter;

ARCHITECTURE a OF Counter IS

	SIGNAL count : unsigned(19 DOWNTO 0) := "00000000000000000000";

BEGIN

	PROCESS(CLK, ASYNCCLRN)
	BEGIN
		IF (ASYNCCLRN = '0') THEN
			count <= "00000000000000000000";
		ELSIF (CLK' EVENT) AND (CLK = '1') THEN
			IF (SYNCCLRN = '0') THEN
				count <= "00000000000000000000";
			ELSE
				count <= count + "1";
			END IF;
		END IF;
	END PROCESS;
	
	Q <= STD_LOGIC_VECTOR(count);

END a;
